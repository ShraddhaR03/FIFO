package fifo_pkg;

`include "uvm_macros.svh" 
import uvm_pkg::*;

`include "seq_item.sv"
`include "op_monitor.sv"
`include "ip_monitor.sv"
`include "ip_driver.sv"
`include "ip_seqr.sv" 
`include "op_agent.sv"
`include "ip_agent.sv"
`include "scoreboard.sv"
`include "coverage_collector.sv"
`include "vseqr.sv"
`include "env.sv"
 `include "seq.sv"
`include "vseq.sv"
 `include "test.sv"

endpackage
